library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity introduction is 
	Port ( switch_0: in STD_LOGIC;
			 switch_1 : in STD_LOGIC;
			 LED_0 : out STD_LOGIC;
			 LED_1 : out STD_LOGIC);
end introduction;

architecture Behavioral of introduction is 
	begin
end Behavioral;
